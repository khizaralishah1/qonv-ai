module store_image();

    reg [7:0] loaded_img [95:0];

endmodule